module top_module( output zero );

// Insert your code here
    assign zero = 0;

endmodule
