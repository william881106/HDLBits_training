module top_module ( input a, input b, output out );
    mod_a U0(a,b,out);
endmodule
